// テストベンチ
// Mux8Way16
module Mux8Way16_tb();
	reg clk = 0;
	reg[15:0] a, b, c, d, e, f, g, h;
	reg[2:0] sel;
	reg[15:0] out;

	parameter RATE = 1;

	always #1 clk = !clk;

	Mux8Way16 mux8Way16(
		.a(a),
		.b(b),
		.c(c),
		.d(d),
		.e(e),
		.f(f),
		.g(g),
		.h(h),
		.sel(sel),
		.out(out)
	);

	initial begin
		$display("start test");
		clk <= 1;

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b000;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b001;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b010;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b011;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b100;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b101;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b110;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0000000000000000; b <= 16'b0000000000000000; c <= 16'b0000000000000000; d <= 16'b0000000000000000; e <= 16'b0000000000000000; f <= 16'b0000000000000000; g <= 16'b0000000000000000; h <= 16'b0000000000000000; sel <= 3'b111;
		#(RATE)
		if (out != 16'b0000000000000000) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b000;
		#(RATE)
		if (out != 16'b0001001000110100) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b001;
		#(RATE)
		if (out != 16'b0010001101000101) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b010;
		#(RATE)
		if (out != 16'b0011010001010110) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b011;
		#(RATE)
		if (out != 16'b0100010101100111) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b100;
		#(RATE)
		if (out != 16'b0101011001111000) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b101;
		#(RATE)
		if (out != 16'b0110011110001001) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b110;
		#(RATE)
		if (out != 16'b0111100010011010) $display("#1 ng");

		#(RATE)
		a <= 16'b0001001000110100; b <= 16'b0010001101000101; c <= 16'b0011010001010110; d <= 16'b0100010101100111; e <= 16'b0101011001111000; f <= 16'b0110011110001001; g <= 16'b0111100010011010; h <= 16'b1000100110101011; sel <= 3'b111;
		#(RATE)
		if (out != 16'b1000100110101011) $display("#1 ng");

		#99999
		$display("success!");
		$stop;
	end

endmodule
