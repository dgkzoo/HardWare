// トップレベル
module HardWare(input clk);
    always @(posedge clk) begin
    end
endmodule
